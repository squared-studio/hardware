// Description
// Author : Foez Ahmed (foez.official@gmail.com)
// This file is part of squared-studio : hardware
// Copyright (c) 2026 squared-studio
// Licensed under the MIT License
// See LICENSE file in the repository root for full license information

module pll_tb;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  localparam int RefDivWidth = 8;
  localparam int FbDivWidth = 12;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////


  logic                   arst_ni;
  logic                   clk_ref_i;
  logic [RefDivWidth-1:0] ref_div_i;
  logic [ FbDivWidth-1:0] fb_div_i;
  logic                   clk_o;
  logic                   locked_o;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INTERFACES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-CLASSES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  pll #(
      .REF_DEV_WIDTH(RefDivWidth),
      .FB_DIV_WIDTH (FbDivWidth)
  ) u_dut (
      .arst_ni  (arst_ni),
      .clk_ref_i(clk_ref_i),
      .ref_div_i(ref_div_i),
      .fb_div_i (fb_div_i),
      .clk_o    (clk_o),
      .locked_o (locked_o)
  );

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  task static apply_reset();
    #100ns;
    arst_ni   <= 0;
    clk_ref_i <= 0;
    ref_div_i <= 0;
    fb_div_i  <= 0;
    #100ns;
    arst_ni <= 1;
    #100ns;
  endtask

  task static start_clock();
    fork
      forever begin
        clk_ref_i <= 1;
        #5ns;
        clk_ref_i <= 0;
        #5ns;
      end
    join_none
    @(posedge clk_ref_i);
  endtask

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin  // main initial

    $dumpfile("pll_tb.vcd");
    $dumpvars(0, pll_tb);

    apply_reset();
    start_clock();

    #10us;

    ref_div_i <= 'd2;

    #10us;

    fb_div_i <= 'd4;

    #10us;

    ref_div_i <= 'd8;
    fb_div_i  <= 'd400;

    #20us;

    $finish;

  end

endmodule
