// Description: This module implements an 8b/10b encoder as per the 8b/10b encoding scheme. It takes
// an 8-bit data input, a control character indicator, and the current running disparity, and
// outputs a 10-bit encoded data, a legality indicator, and the updated running disparity.
// -------------------------------------------------------------------------------------------------
// Author : Foez Ahmed (foez.official@gmail.com)
// This file is part of squared-studio : hardware
// Copyright (c) 2026 squared-studio
// Licensed under the MIT License
// See LICENSE file in the repository root for full license information


module encoder_8b10b (
    // 8-bit input data to be encoded
    input logic [7:0] data_i,
    // Control character indicator (1 for K-character, 0 for D-character)
    input logic k_char_i,
    // Current running disparity (0 for RD-, 1 for RD+)
    input logic running_disparity_i,

    // 10-bit encoded output data
    output logic [9:0] data_o,
    // Indicates if the input combination is legal (1 for legal, 0 for illegal)
    output logic       is_legal_o,
    // Updated running disparity after encoding (0 for RD-, 1 for RD+)
    output logic       running_disparity_o
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // Combinational logic block for 8b/10b encoding
  // The 'always_comb' block infers combinational logic, meaning outputs react immediately to input changes.
  always_comb begin
    case ({
      data_i, k_char_i, running_disparity_i
    })
      10'b00000000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001110100_1_1;  // D00.0 -
      10'b00000000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110001011_1_0;  // D00.0 +
      10'b00000001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111010100_1_1;  // D01.0 -
      10'b00000001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000101011_1_0;  // D01.0 +
      10'b00000010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011010100_1_1;  // D02.0 -
      10'b00000010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100101011_1_0;  // D02.0 +
      10'b00000011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100011011_1_1;  // D03.0 -
      10'b00000011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100010100_1_0;  // D03.0 +
      10'b00000100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101010100_1_1;  // D04.0 -
      10'b00000100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010101011_1_0;  // D04.0 +
      10'b00000101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010011011_1_1;  // D05.0 -
      10'b00000101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010010100_1_0;  // D05.0 +
      10'b00000110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110011011_1_1;  // D06.0 -
      10'b00000110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110010100_1_0;  // D06.0 +
      10'b00000111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110001011_1_1;  // D07.0 -
      10'b00000111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001110100_1_0;  // D07.0 +
      10'b00001000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110010100_1_1;  // D08.0 -
      10'b00001000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001101011_1_0;  // D08.0 +
      10'b00001001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001011011_1_1;  // D09.0 -
      10'b00001001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001010100_1_0;  // D09.0 +
      10'b00001010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101011011_1_1;  // D10.0 -
      10'b00001010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101010100_1_0;  // D10.0 +
      10'b00001011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101001011_1_1;  // D11.0 -
      10'b00001011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1101000100_1_0;  // D11.0 +
      10'b00001100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011011011_1_1;  // D12.0 -
      10'b00001100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011010100_1_0;  // D12.0 +
      10'b00001101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011001011_1_1;  // D13.0 -
      10'b00001101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1011000100_1_0;  // D13.0 +
      10'b00001110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111001011_1_1;  // D14.0 -
      10'b00001110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0111000100_1_0;  // D14.0 +
      10'b00001111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101110100_1_1;  // D15.0 -
      10'b00001111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010001011_1_0;  // D15.0 +
      10'b00010000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110110100_1_1;  // D16.0 -
      10'b00010000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001001011_1_0;  // D16.0 +
      10'b00010001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1000111011_1_1;  // D17.0 -
      10'b00010001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000110100_1_0;  // D17.0 +
      10'b00010010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0100111011_1_1;  // D18.0 -
      10'b00010010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100110100_1_0;  // D18.0 +
      10'b00010011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100101011_1_1;  // D19.0 -
      10'b00010011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100100100_1_0;  // D19.0 +
      10'b00010100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0010111011_1_1;  // D20.0 -
      10'b00010100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010110100_1_0;  // D20.0 +
      10'b00010101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010101011_1_1;  // D21.0 -
      10'b00010101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010100100_1_0;  // D21.0 +
      10'b00010110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110101011_1_1;  // D22.0 -
      10'b00010110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110100100_1_0;  // D22.0 +
      10'b00010111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110100100_1_1;  // D23.0 -
      10'b00010111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001011011_1_0;  // D23.0 +
      10'b00011000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100110100_1_1;  // D24.0 -
      10'b00011000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011001011_1_0;  // D24.0 +
      10'b00011001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001101011_1_1;  // D25.0 -
      10'b00011001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001100100_1_0;  // D25.0 +
      10'b00011010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101101011_1_1;  // D26.0 -
      10'b00011010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101100100_1_0;  // D26.0 +
      10'b00011011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101100100_1_1;  // D27.0 -
      10'b00011011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010011011_1_0;  // D27.0 +
      10'b00011100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011101011_1_1;  // D28.0 -
      10'b00011100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011100100_1_0;  // D28.0 +
      10'b00011101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011100100_1_1;  // D29.0 -
      10'b00011101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100011011_1_0;  // D29.0 +
      10'b00011110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111100100_1_1;  // D30.0 -
      10'b00011110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000011011_1_0;  // D30.0 +
      10'b00011111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010110100_1_1;  // D31.0 -
      10'b00011111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101001011_1_0;  // D31.0 +
      10'b00100000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001111001_1_1;  // D00.1 -
      10'b00100000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110001001_1_0;  // D00.1 +
      10'b00100001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111011001_1_1;  // D01.1 -
      10'b00100001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000101001_1_0;  // D01.1 +
      10'b00100010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011011001_1_1;  // D02.1 -
      10'b00100010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100101001_1_0;  // D02.1 +
      10'b00100011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100011001_1_0;  // D03.1 +
      10'b00100011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100011001_1_1;  // D03.1 -
      10'b00100100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101011001_1_1;  // D04.1 -
      10'b00100100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010101001_1_0;  // D04.1 +
      10'b00100101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010011001_1_0;  // D05.1 +
      10'b00100101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010011001_1_1;  // D05.1 -
      10'b00100110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110011001_1_0;  // D06.1 +
      10'b00100110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110011001_1_1;  // D06.1 -
      10'b00100111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110001001_1_1;  // D07.1 -
      10'b00100111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001111001_1_0;  // D07.1 +
      10'b00101000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110011001_1_1;  // D08.1 -
      10'b00101000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001101001_1_0;  // D08.1 +
      10'b00101001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001011001_1_0;  // D09.1 +
      10'b00101001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001011001_1_1;  // D09.1 -
      10'b00101010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101011001_1_0;  // D10.1 +
      10'b00101010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101011001_1_1;  // D10.1 -
      10'b00101011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101001001_1_0;  // D11.1 +
      10'b00101011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1101001001_1_1;  // D11.1 -
      10'b00101100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011011001_1_0;  // D12.1 +
      10'b00101100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011011001_1_1;  // D12.1 -
      10'b00101101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011001001_1_0;  // D13.1 +
      10'b00101101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1011001001_1_1;  // D13.1 -
      10'b00101110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111001001_1_0;  // D14.1 +
      10'b00101110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0111001001_1_1;  // D14.1 -
      10'b00101111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101111001_1_1;  // D15.1 -
      10'b00101111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010001001_1_0;  // D15.1 +
      10'b00110000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110111001_1_1;  // D16.1 -
      10'b00110000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001001001_1_0;  // D16.1 +
      10'b00110001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1000111001_1_0;  // D17.1 +
      10'b00110001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000111001_1_1;  // D17.1 -
      10'b00110010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0100111001_1_0;  // D18.1 +
      10'b00110010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100111001_1_1;  // D18.1 -
      10'b00110011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100101001_1_0;  // D19.1 +
      10'b00110011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100101001_1_1;  // D19.1 -
      10'b00110100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0010111001_1_0;  // D20.1 +
      10'b00110100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010111001_1_1;  // D20.1 -
      10'b00110101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010101001_1_0;  // D21.1 +
      10'b00110101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010101001_1_1;  // D21.1 -
      10'b00110110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110101001_1_0;  // D22.1 +
      10'b00110110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110101001_1_1;  // D22.1 -
      10'b00110111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110101001_1_1;  // D23.1 -
      10'b00110111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001011001_1_0;  // D23.1 +
      10'b00111000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100111001_1_1;  // D24.1 -
      10'b00111000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011001001_1_0;  // D24.1 +
      10'b00111001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001101001_1_0;  // D25.1 +
      10'b00111001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001101001_1_1;  // D25.1 -
      10'b00111010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101101001_1_0;  // D26.1 +
      10'b00111010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101101001_1_1;  // D26.1 -
      10'b00111011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101101001_1_1;  // D27.1 -
      10'b00111011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010011001_1_0;  // D27.1 +
      10'b00111100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011101001_1_0;  // D28.1 +
      10'b00111100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011101001_1_1;  // D28.1 -
      10'b00111101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011101001_1_1;  // D29.1 -
      10'b00111101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100011001_1_0;  // D29.1 +
      10'b00111110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111101001_1_1;  // D30.1 -
      10'b00111110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000011001_1_0;  // D30.1 +
      10'b00111111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010111001_1_1;  // D31.1 -
      10'b00111111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101001001_1_0;  // D31.1 +
      10'b01000000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001110101_1_1;  // D00.2 -
      10'b01000000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110000101_1_0;  // D00.2 +
      10'b01000001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111010101_1_1;  // D01.2 -
      10'b01000001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000100101_1_0;  // D01.2 +
      10'b01000010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011010101_1_1;  // D02.2 -
      10'b01000010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100100101_1_0;  // D02.2 +
      10'b01000011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100010101_1_0;  // D03.2 +
      10'b01000011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100010101_1_1;  // D03.2 -
      10'b01000100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101010101_1_1;  // D04.2 -
      10'b01000100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010100101_1_0;  // D04.2 +
      10'b01000101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010010101_1_0;  // D05.2 +
      10'b01000101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010010101_1_1;  // D05.2 -
      10'b01000110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110010101_1_0;  // D06.2 +
      10'b01000110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110010101_1_1;  // D06.2 -
      10'b01000111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110000101_1_1;  // D07.2 -
      10'b01000111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001110101_1_0;  // D07.2 +
      10'b01001000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110010101_1_1;  // D08.2 -
      10'b01001000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001100101_1_0;  // D08.2 +
      10'b01001001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001010101_1_0;  // D09.2 +
      10'b01001001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001010101_1_1;  // D09.2 -
      10'b01001010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101010101_1_0;  // D10.2 +
      10'b01001010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101010101_1_1;  // D10.2 -
      10'b01001011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101000101_1_0;  // D11.2 +
      10'b01001011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1101000101_1_1;  // D11.2 -
      10'b01001100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011010101_1_0;  // D12.2 +
      10'b01001100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011010101_1_1;  // D12.2 -
      10'b01001101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011000101_1_0;  // D13.2 +
      10'b01001101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1011000101_1_1;  // D13.2 -
      10'b01001110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111000101_1_0;  // D14.2 +
      10'b01001110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0111000101_1_1;  // D14.2 -
      10'b01001111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101110101_1_1;  // D15.2 -
      10'b01001111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010000101_1_0;  // D15.2 +
      10'b01010000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110110101_1_1;  // D16.2 -
      10'b01010000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001000101_1_0;  // D16.2 +
      10'b01010001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1000110101_1_0;  // D17.2 +
      10'b01010001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000110101_1_1;  // D17.2 -
      10'b01010010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0100110101_1_0;  // D18.2 +
      10'b01010010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100110101_1_1;  // D18.2 -
      10'b01010011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100100101_1_0;  // D19.2 +
      10'b01010011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100100101_1_1;  // D19.2 -
      10'b01010100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0010110101_1_0;  // D20.2 +
      10'b01010100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010110101_1_1;  // D20.2 -
      10'b01010101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010100101_1_0;  // D21.2 +
      10'b01010101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010100101_1_1;  // D21.2 -
      10'b01010110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110100101_1_0;  // D22.2 +
      10'b01010110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110100101_1_1;  // D22.2 -
      10'b01010111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110100101_1_1;  // D23.2 -
      10'b01010111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001010101_1_0;  // D23.2 +
      10'b01011000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100110101_1_1;  // D24.2 -
      10'b01011000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011000101_1_0;  // D24.2 +
      10'b01011001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001100101_1_0;  // D25.2 +
      10'b01011001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001100101_1_1;  // D25.2 -
      10'b01011010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101100101_1_0;  // D26.2 +
      10'b01011010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101100101_1_1;  // D26.2 -
      10'b01011011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101100101_1_1;  // D27.2 -
      10'b01011011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010010101_1_0;  // D27.2 +
      10'b01011100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011100101_1_0;  // D28.2 +
      10'b01011100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011100101_1_1;  // D28.2 -
      10'b01011101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011100101_1_1;  // D29.2 -
      10'b01011101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100010101_1_0;  // D29.2 +
      10'b01011110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111100101_1_1;  // D30.2 -
      10'b01011110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000010101_1_0;  // D30.2 +
      10'b01011111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010110101_1_1;  // D31.2 -
      10'b01011111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101000101_1_0;  // D31.2 +
      10'b01100000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001110011_1_1;  // D00.3 -
      10'b01100000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110001100_1_0;  // D00.3 +
      10'b01100001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111010011_1_1;  // D01.3 -
      10'b01100001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000101100_1_0;  // D01.3 +
      10'b01100010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011010011_1_1;  // D02.3 -
      10'b01100010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100101100_1_0;  // D02.3 +
      10'b01100011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100011100_1_1;  // D03.3 -
      10'b01100011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100010011_1_0;  // D03.3 +
      10'b01100100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101010011_1_1;  // D04.3 -
      10'b01100100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010101100_1_0;  // D04.3 +
      10'b01100101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010011100_1_1;  // D05.3 -
      10'b01100101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010010011_1_0;  // D05.3 +
      10'b01100110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110011100_1_1;  // D06.3 -
      10'b01100110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110010011_1_0;  // D06.3 +
      10'b01100111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110001100_1_1;  // D07.3 -
      10'b01100111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001110011_1_0;  // D07.3 +
      10'b01101000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110010011_1_1;  // D08.3 -
      10'b01101000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001101100_1_0;  // D08.3 +
      10'b01101001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001011100_1_1;  // D09.3 -
      10'b01101001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001010011_1_0;  // D09.3 +
      10'b01101010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101011100_1_1;  // D10.3 -
      10'b01101010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101010011_1_0;  // D10.3 +
      10'b01101011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101001100_1_1;  // D11.3 -
      10'b01101011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1101000011_1_0;  // D11.3 +
      10'b01101100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011011100_1_1;  // D12.3 -
      10'b01101100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011010011_1_0;  // D12.3 +
      10'b01101101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011001100_1_1;  // D13.3 -
      10'b01101101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1011000011_1_0;  // D13.3 +
      10'b01101110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111001100_1_1;  // D14.3 -
      10'b01101110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0111000011_1_0;  // D14.3 +
      10'b01101111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101110011_1_1;  // D15.3 -
      10'b01101111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010001100_1_0;  // D15.3 +
      10'b01110000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110110011_1_1;  // D16.3 -
      10'b01110000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001001100_1_0;  // D16.3 +
      10'b01110001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1000111100_1_1;  // D17.3 -
      10'b01110001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000110011_1_0;  // D17.3 +
      10'b01110010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0100111100_1_1;  // D18.3 -
      10'b01110010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100110011_1_0;  // D18.3 +
      10'b01110011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100101100_1_1;  // D19.3 -
      10'b01110011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100100011_1_0;  // D19.3 +
      10'b01110100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0010111100_1_1;  // D20.3 -
      10'b01110100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010110011_1_0;  // D20.3 +
      10'b01110101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010101100_1_1;  // D21.3 -
      10'b01110101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010100011_1_0;  // D21.3 +
      10'b01110110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110101100_1_1;  // D22.3 -
      10'b01110110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110100011_1_0;  // D22.3 +
      10'b01110111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110100011_1_1;  // D23.3 -
      10'b01110111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001011100_1_0;  // D23.3 +
      10'b01111000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100110011_1_1;  // D24.3 -
      10'b01111000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011001100_1_0;  // D24.3 +
      10'b01111001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001101100_1_1;  // D25.3 -
      10'b01111001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001100011_1_0;  // D25.3 +
      10'b01111010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101101100_1_1;  // D26.3 -
      10'b01111010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101100011_1_0;  // D26.3 +
      10'b01111011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101100011_1_1;  // D27.3 -
      10'b01111011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010011100_1_0;  // D27.3 +
      10'b01111100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011101100_1_1;  // D28.3 -
      10'b01111100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011100011_1_0;  // D28.3 +
      10'b01111101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011100011_1_1;  // D29.3 -
      10'b01111101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100011100_1_0;  // D29.3 +
      10'b01111110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111100011_1_1;  // D30.3 -
      10'b01111110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000011100_1_0;  // D30.3 +
      10'b01111111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010110011_1_1;  // D31.3 -
      10'b01111111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101001100_1_0;  // D31.3 +
      10'b10000000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001110010_1_1;  // D00.4 -
      10'b10000000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110001101_1_0;  // D00.4 +
      10'b10000001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111010010_1_1;  // D01.4 -
      10'b10000001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000101101_1_0;  // D01.4 +
      10'b10000010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011010010_1_1;  // D02.4 -
      10'b10000010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100101101_1_0;  // D02.4 +
      10'b10000011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100011101_1_1;  // D03.4 -
      10'b10000011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100010010_1_0;  // D03.4 +
      10'b10000100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101010010_1_1;  // D04.4 -
      10'b10000100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010101101_1_0;  // D04.4 +
      10'b10000101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010011101_1_1;  // D05.4 -
      10'b10000101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010010010_1_0;  // D05.4 +
      10'b10000110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110011101_1_1;  // D06.4 -
      10'b10000110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110010010_1_0;  // D06.4 +
      10'b10000111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110001101_1_1;  // D07.4 -
      10'b10000111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001110010_1_0;  // D07.4 +
      10'b10001000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110010010_1_1;  // D08.4 -
      10'b10001000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001101101_1_0;  // D08.4 +
      10'b10001001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001011101_1_1;  // D09.4 -
      10'b10001001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001010010_1_0;  // D09.4 +
      10'b10001010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101011101_1_1;  // D10.4 -
      10'b10001010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101010010_1_0;  // D10.4 +
      10'b10001011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101001101_1_1;  // D11.4 -
      10'b10001011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1101000010_1_0;  // D11.4 +
      10'b10001100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011011101_1_1;  // D12.4 -
      10'b10001100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011010010_1_0;  // D12.4 +
      10'b10001101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011001101_1_1;  // D13.4 -
      10'b10001101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1011000010_1_0;  // D13.4 +
      10'b10001110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111001101_1_1;  // D14.4 -
      10'b10001110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0111000010_1_0;  // D14.4 +
      10'b10001111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101110010_1_1;  // D15.4 -
      10'b10001111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010001101_1_0;  // D15.4 +
      10'b10010000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110110010_1_1;  // D16.4 -
      10'b10010000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001001101_1_0;  // D16.4 +
      10'b10010001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1000111101_1_1;  // D17.4 -
      10'b10010001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000110010_1_0;  // D17.4 +
      10'b10010010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0100111101_1_1;  // D18.4 -
      10'b10010010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100110010_1_0;  // D18.4 +
      10'b10010011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100101101_1_1;  // D19.4 -
      10'b10010011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100100010_1_0;  // D19.4 +
      10'b10010100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0010111101_1_1;  // D20.4 -
      10'b10010100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010110010_1_0;  // D20.4 +
      10'b10010101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010101101_1_1;  // D21.4 -
      10'b10010101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010100010_1_0;  // D21.4 +
      10'b10010110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110101101_1_1;  // D22.4 -
      10'b10010110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110100010_1_0;  // D22.4 +
      10'b10010111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110100010_1_1;  // D23.4 -
      10'b10010111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001011101_1_0;  // D23.4 +
      10'b10011000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100110010_1_1;  // D24.4 -
      10'b10011000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011001101_1_0;  // D24.4 +
      10'b10011001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001101101_1_1;  // D25.4 -
      10'b10011001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001100010_1_0;  // D25.4 +
      10'b10011010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101101101_1_1;  // D26.4 -
      10'b10011010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101100010_1_0;  // D26.4 +
      10'b10011011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101100010_1_1;  // D27.4 -
      10'b10011011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010011101_1_0;  // D27.4 +
      10'b10011100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011101101_1_1;  // D28.4 -
      10'b10011100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011100010_1_0;  // D28.4 +
      10'b10011101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011100010_1_1;  // D29.4 -
      10'b10011101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100011101_1_0;  // D29.4 +
      10'b10011110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111100010_1_1;  // D30.4 -
      10'b10011110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000011101_1_0;  // D30.4 +
      10'b10011111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010110010_1_1;  // D31.4 -
      10'b10011111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101001101_1_0;  // D31.4 +
      10'b10100000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001111010_1_1;  // D00.5 -
      10'b10100000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110001010_1_0;  // D00.5 +
      10'b10100001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111011010_1_1;  // D01.5 -
      10'b10100001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000101010_1_0;  // D01.5 +
      10'b10100010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011011010_1_1;  // D02.5 -
      10'b10100010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100101010_1_0;  // D02.5 +
      10'b10100011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100011010_1_0;  // D03.5 +
      10'b10100011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100011010_1_1;  // D03.5 -
      10'b10100100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101011010_1_1;  // D04.5 -
      10'b10100100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010101010_1_0;  // D04.5 +
      10'b10100101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010011010_1_0;  // D05.5 +
      10'b10100101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010011010_1_1;  // D05.5 -
      10'b10100110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110011010_1_0;  // D06.5 +
      10'b10100110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110011010_1_1;  // D06.5 -
      10'b10100111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110001010_1_1;  // D07.5 -
      10'b10100111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001111010_1_0;  // D07.5 +
      10'b10101000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110011010_1_1;  // D08.5 -
      10'b10101000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001101010_1_0;  // D08.5 +
      10'b10101001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001011010_1_0;  // D09.5 +
      10'b10101001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001011010_1_1;  // D09.5 -
      10'b10101010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101011010_1_0;  // D10.5 +
      10'b10101010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101011010_1_1;  // D10.5 -
      10'b10101011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101001010_1_0;  // D11.5 +
      10'b10101011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1101001010_1_1;  // D11.5 -
      10'b10101100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011011010_1_0;  // D12.5 +
      10'b10101100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011011010_1_1;  // D12.5 -
      10'b10101101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011001010_1_0;  // D13.5 +
      10'b10101101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1011001010_1_1;  // D13.5 -
      10'b10101110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111001010_1_0;  // D14.5 +
      10'b10101110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0111001010_1_1;  // D14.5 -
      10'b10101111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101111010_1_1;  // D15.5 -
      10'b10101111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010001010_1_0;  // D15.5 +
      10'b10110000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110111010_1_1;  // D16.5 -
      10'b10110000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001001010_1_0;  // D16.5 +
      10'b10110001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1000111010_1_0;  // D17.5 +
      10'b10110001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000111010_1_1;  // D17.5 -
      10'b10110010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0100111010_1_0;  // D18.5 +
      10'b10110010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100111010_1_1;  // D18.5 -
      10'b10110011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100101010_1_0;  // D19.5 +
      10'b10110011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100101010_1_1;  // D19.5 -
      10'b10110100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0010111010_1_0;  // D20.5 +
      10'b10110100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010111010_1_1;  // D20.5 -
      10'b10110101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010101010_1_0;  // D21.5 +
      10'b10110101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010101010_1_1;  // D21.5 -
      10'b10110110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110101010_1_0;  // D22.5 +
      10'b10110110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110101010_1_1;  // D22.5 -
      10'b10110111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110101010_1_1;  // D23.5 -
      10'b10110111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001011010_1_0;  // D23.5 +
      10'b10111000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100111010_1_1;  // D24.5 -
      10'b10111000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011001010_1_0;  // D24.5 +
      10'b10111001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001101010_1_0;  // D25.5 +
      10'b10111001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001101010_1_1;  // D25.5 -
      10'b10111010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101101010_1_0;  // D26.5 +
      10'b10111010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101101010_1_1;  // D26.5 -
      10'b10111011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101101010_1_1;  // D27.5 -
      10'b10111011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010011010_1_0;  // D27.5 +
      10'b10111100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011101010_1_0;  // D28.5 +
      10'b10111100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011101010_1_1;  // D28.5 -
      10'b10111101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011101010_1_1;  // D29.5 -
      10'b10111101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100011010_1_0;  // D29.5 +
      10'b10111110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111101010_1_1;  // D30.5 -
      10'b10111110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000011010_1_0;  // D30.5 +
      10'b10111111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010111010_1_1;  // D31.5 -
      10'b10111111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101001010_1_0;  // D31.5 +
      10'b11000000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001110110_1_1;  // D00.6 -
      10'b11000000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110000110_1_0;  // D00.6 +
      10'b11000001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111010110_1_1;  // D01.6 -
      10'b11000001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000100110_1_0;  // D01.6 +
      10'b11000010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011010110_1_1;  // D02.6 -
      10'b11000010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100100110_1_0;  // D02.6 +
      10'b11000011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100010110_1_0;  // D03.6 +
      10'b11000011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100010110_1_1;  // D03.6 -
      10'b11000100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101010110_1_1;  // D04.6 -
      10'b11000100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010100110_1_0;  // D04.6 +
      10'b11000101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010010110_1_0;  // D05.6 +
      10'b11000101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010010110_1_1;  // D05.6 -
      10'b11000110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110010110_1_0;  // D06.6 +
      10'b11000110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110010110_1_1;  // D06.6 -
      10'b11000111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110000110_1_1;  // D07.6 -
      10'b11000111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001110110_1_0;  // D07.6 +
      10'b11001000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110010110_1_1;  // D08.6 -
      10'b11001000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001100110_1_0;  // D08.6 +
      10'b11001001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001010110_1_0;  // D09.6 +
      10'b11001001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001010110_1_1;  // D09.6 -
      10'b11001010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101010110_1_0;  // D10.6 +
      10'b11001010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101010110_1_1;  // D10.6 -
      10'b11001011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101000110_1_0;  // D11.6 +
      10'b11001011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1101000110_1_1;  // D11.6 -
      10'b11001100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011010110_1_0;  // D12.6 +
      10'b11001100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011010110_1_1;  // D12.6 -
      10'b11001101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011000110_1_0;  // D13.6 +
      10'b11001101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1011000110_1_1;  // D13.6 -
      10'b11001110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111000110_1_0;  // D14.6 +
      10'b11001110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0111000110_1_1;  // D14.6 -
      10'b11001111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101110110_1_1;  // D15.6 -
      10'b11001111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010000110_1_0;  // D15.6 +
      10'b11010000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110110110_1_1;  // D16.6 -
      10'b11010000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001000110_1_0;  // D16.6 +
      10'b11010001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1000110110_1_0;  // D17.6 +
      10'b11010001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000110110_1_1;  // D17.6 -
      10'b11010010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0100110110_1_0;  // D18.6 +
      10'b11010010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100110110_1_1;  // D18.6 -
      10'b11010011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100100110_1_0;  // D19.6 +
      10'b11010011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100100110_1_1;  // D19.6 -
      10'b11010100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0010110110_1_0;  // D20.6 +
      10'b11010100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010110110_1_1;  // D20.6 -
      10'b11010101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010100110_1_0;  // D21.6 +
      10'b11010101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010100110_1_1;  // D21.6 -
      10'b11010110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110100110_1_0;  // D22.6 +
      10'b11010110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110100110_1_1;  // D22.6 -
      10'b11010111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110100110_1_1;  // D23.6 -
      10'b11010111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001010110_1_0;  // D23.6 +
      10'b11011000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100110110_1_1;  // D24.6 -
      10'b11011000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011000110_1_0;  // D24.6 +
      10'b11011001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001100110_1_0;  // D25.6 +
      10'b11011001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001100110_1_1;  // D25.6 -
      10'b11011010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101100110_1_0;  // D26.6 +
      10'b11011010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101100110_1_1;  // D26.6 -
      10'b11011011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101100110_1_1;  // D27.6 -
      10'b11011011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010010110_1_0;  // D27.6 +
      10'b11011100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011100110_1_0;  // D28.6 +
      10'b11011100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011100110_1_1;  // D28.6 -
      10'b11011101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011100110_1_1;  // D29.6 -
      10'b11011101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100010110_1_0;  // D29.6 +
      10'b11011110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111100110_1_1;  // D30.6 -
      10'b11011110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000010110_1_0;  // D30.6 +
      10'b11011111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010110110_1_1;  // D31.6 -
      10'b11011111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101000110_1_0;  // D31.6 +
      10'b11100000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001110001_1_1;  // D00.7 -
      10'b11100000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110001110_1_0;  // D00.7 +
      10'b11100001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111010001_1_1;  // D01.7 -
      10'b11100001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000101110_1_0;  // D01.7 +
      10'b11100010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011010001_1_1;  // D02.7 -
      10'b11100010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100101110_1_0;  // D02.7 +
      10'b11100011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100011110_1_1;  // D03.7 -
      10'b11100011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100010001_1_0;  // D03.7 +
      10'b11100100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101010001_1_1;  // D04.7 -
      10'b11100100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010101110_1_0;  // D04.7 +
      10'b11100101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010011110_1_1;  // D05.7 -
      10'b11100101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010010001_1_0;  // D05.7 +
      10'b11100110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110011110_1_1;  // D06.7 -
      10'b11100110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110010001_1_0;  // D06.7 +
      10'b11100111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110001110_1_1;  // D07.7 -
      10'b11100111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001110001_1_0;  // D07.7 +
      10'b11101000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110010001_1_1;  // D08.7 -
      10'b11101000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001101110_1_0;  // D08.7 +
      10'b11101001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001011110_1_1;  // D09.7 -
      10'b11101001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001010001_1_0;  // D09.7 +
      10'b11101010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101011110_1_1;  // D10.7 -
      10'b11101010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101010001_1_0;  // D10.7 +
      10'b11101011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101001110_1_1;  // D11.7 -
      10'b11101011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1101001000_1_0;  // D11.7 +
      10'b11101100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011011110_1_1;  // D12.7 -
      10'b11101100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011010001_1_0;  // D12.7 +
      10'b11101101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011001110_1_1;  // D13.7 -
      10'b11101101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1011001000_1_0;  // D13.7 +
      10'b11101110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111001110_1_1;  // D14.7 -
      10'b11101110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0111001000_1_0;  // D14.7 +
      10'b11101111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101110001_1_1;  // D15.7 -
      10'b11101111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010001110_1_0;  // D15.7 +
      10'b11110000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110110001_1_1;  // D16.7 -
      10'b11110000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001001110_1_0;  // D16.7 +
      10'b11110001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1000110111_1_1;  // D17.7 -
      10'b11110001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000110001_1_0;  // D17.7 +
      10'b11110010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0100110111_1_1;  // D18.7 -
      10'b11110010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100110001_1_0;  // D18.7 +
      10'b11110011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100101110_1_1;  // D19.7 -
      10'b11110011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100100001_1_0;  // D19.7 +
      10'b11110100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0010110111_1_1;  // D20.7 -
      10'b11110100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010110001_1_0;  // D20.7 +
      10'b11110101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010101110_1_1;  // D21.7 -
      10'b11110101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1010100001_1_0;  // D21.7 +
      10'b11110110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0110101110_1_1;  // D22.7 -
      10'b11110110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0110100001_1_0;  // D22.7 +
      10'b11110111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110100001_1_1;  // D23.7 -
      10'b11110111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001011110_1_0;  // D23.7 +
      10'b11111000_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1100110001_1_1;  // D24.7 -
      10'b11111000_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011001110_1_0;  // D24.7 +
      10'b11111001_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1001101110_1_1;  // D25.7 -
      10'b11111001_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1001100001_1_0;  // D25.7 +
      10'b11111010_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0101101110_1_1;  // D26.7 -
      10'b11111010_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101100001_1_0;  // D26.7 +
      10'b11111011_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101100001_1_1;  // D27.7 -
      10'b11111011_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010011110_1_0;  // D27.7 +
      10'b11111100_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011101110_1_1;  // D28.7 -
      10'b11111100_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0011100001_1_0;  // D28.7 +
      10'b11111101_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011100001_1_1;  // D29.7 -
      10'b11111101_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100011110_1_0;  // D29.7 +
      10'b11111110_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111100001_1_1;  // D30.7 -
      10'b11111110_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000011110_1_0;  // D30.7 +
      10'b11111111_0_0: {data_o, is_legal_o, running_disparity_o} = 12'b1010110001_1_1;  // D31.7 -
      10'b11111111_0_1: {data_o, is_legal_o, running_disparity_o} = 12'b0101001110_1_0;  // D31.7 +
      10'b00011100_1_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011110100_1_1;  // K28.0 -
      10'b00011100_1_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100001011_1_0;  // K28.0 +
      10'b00111100_1_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011111001_1_1;  // K28.1 -
      10'b00111100_1_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100000110_1_0;  // K28.1 +
      10'b01011100_1_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011110101_1_1;  // K28.2 -
      10'b01011100_1_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100001010_1_0;  // K28.2 +
      10'b01111100_1_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011110011_1_1;  // K28.3 -
      10'b01111100_1_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100001100_1_0;  // K28.3 +
      10'b10011100_1_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011110010_1_1;  // K28.4 -
      10'b10011100_1_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100001101_1_0;  // K28.4 +
      10'b10111100_1_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011111010_1_1;  // K28.5 -
      10'b10111100_1_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100000101_1_0;  // K28.5 +
      10'b11011100_1_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011110110_1_1;  // K28.6 -
      10'b11011100_1_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100001001_1_0;  // K28.6 +
      10'b11111100_1_0: {data_o, is_legal_o, running_disparity_o} = 12'b0011111000_1_1;  // K28.7 -
      10'b11111100_1_1: {data_o, is_legal_o, running_disparity_o} = 12'b1100000111_1_0;  // K28.7 +
      10'b11110111_1_0: {data_o, is_legal_o, running_disparity_o} = 12'b1110101000_1_1;  // K23.7 -
      10'b11110111_1_1: {data_o, is_legal_o, running_disparity_o} = 12'b0001010111_1_0;  // K23.7 +
      10'b11111011_1_0: {data_o, is_legal_o, running_disparity_o} = 12'b1101101000_1_1;  // K27.7 -
      10'b11111011_1_1: {data_o, is_legal_o, running_disparity_o} = 12'b0010010111_1_0;  // K27.7 +
      10'b11111101_1_0: {data_o, is_legal_o, running_disparity_o} = 12'b1011101000_1_1;  // K29.7 -
      10'b11111101_1_1: {data_o, is_legal_o, running_disparity_o} = 12'b0100010111_1_0;  // K29.7 +
      10'b11111110_1_0: {data_o, is_legal_o, running_disparity_o} = 12'b0111101000_1_1;  // K30.7 -
      10'b11111110_1_1: {data_o, is_legal_o, running_disparity_o} = 12'b1000010111_1_0;  // K30.7 +
      default:  // ERROR
      {data_o, is_legal_o, running_disparity_o} = {11'b0000000000_0, running_disparity_i};
    endcase
  end

endmodule
