// Description
// Author : Foez Ahmed (foez.official@gmail.com)
// This file is part of squared-studio : hardware
// Copyright (c) 2026 squared-studio
// Licensed under the MIT License
// See LICENSE file in the repository root for full license information

module pll_tb;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  localparam int REF_DEV_WIDTH = 4;
  localparam int FB_DIV_WIDTH = 8;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////


  logic                     arst_ni;
  logic                     clk_ref_i;
  logic [REF_DEV_WIDTH-1:0] refdiv_i;
  logic [ FB_DIV_WIDTH-1:0] fbdiv_i;
  logic                     clk_o;
  logic                     locked_o;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INTERFACES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-CLASSES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  pll #(
      .REF_DEV_WIDTH(REF_DEV_WIDTH),
      .FB_DIV_WIDTH (FB_DIV_WIDTH)
  ) u_dut (
      .arst_ni  (arst_ni),
      .clk_ref_i(clk_ref_i),
      .refdiv_i (refdiv_i),
      .fbdiv_i  (fbdiv_i),
      .clk_o    (clk_o),
      .locked_o (locked_o)
  );

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  task static apply_reset();
    #100ns;
    arst_ni   <= 0;
    clk_ref_i <= 0;
    refdiv_i  <= 0;
    fbdiv_i   <= 0;
    #100ns;
    arst_ni <= 1;
    #100ns;
  endtask

  task static start_clock();
    fork
      forever begin
        clk_ref_i <= 1;
        #5ns;
        clk_ref_i <= 0;
        #5ns;
      end
    join_none
    @(posedge clk_ref_i);
  endtask

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin  // main initial

    $dumpfile("pll_tb.vcd");
    $dumpvars(0, pll_tb);

    apply_reset();
    start_clock();

    #10us;
    
    refdiv_i <= 4'd2;

    #10us;
    
    fbdiv_i <= 8'd4;

    #10us;
    
    refdiv_i <= 4'd8;
    fbdiv_i <= 8'd200;

    #10us;

    $finish;

  end

endmodule
