interface dummy_intf;
  
endinterface
