package dummy_pkg;
  
endpackage
