// Author : Foez Ahmed (foez.official@gmail.com)
// This file is part of squared-studio : hardware
// Copyright (c) 2025 squared-studio
// Licensed under the MIT License
// See LICENSE file in the repository root for full license information

