// Description
// Author : Foez Ahmed (foez.official@gmail.com)
// This file is part of squared-studio : hardware
// Copyright (c) 2026 squared-studio
// Licensed under the MIT License
// See LICENSE file in the repository root for full license information

module pll_tb;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-LOCALPARAMS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  localparam int RefDivWidth = 8;
  localparam int FbDivWidth = 12;

  localparam real RefFreq = 100e6;  // 100 MHz

  localparam real MinOutFreq = 1e6;  // 1 MHz
  localparam real MaxOutFreq = 10e9;  // 10 GHz

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-TYPEDEFS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SIGNALS
  //////////////////////////////////////////////////////////////////////////////////////////////////


  logic                   arst_ni;
  logic                   clk_ref_i;
  logic [RefDivWidth-1:0] ref_div_i;
  logic [ FbDivWidth-1:0] fb_div_i;
  logic                   clk_o;
  logic                   locked_o;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-VARIABLES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  bit                     test_passed;

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-INTERFACES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-CLASSES
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-RTLS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  pll #(
      .REF_DEV_WIDTH(RefDivWidth),
      .FB_DIV_WIDTH (FbDivWidth)
  ) u_dut (
      .arst_ni  (arst_ni),
      .clk_ref_i(clk_ref_i),
      .ref_div_i(ref_div_i),
      .fb_div_i (fb_div_i),
      .clk_o    (clk_o),
      .locked_o (locked_o)
  );

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-METHODS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  task static apply_reset();
    #100ns;
    arst_ni   <= 0;
    clk_ref_i <= 0;
    ref_div_i <= 0;
    fb_div_i  <= 0;
    #100ns;
    arst_ni <= 1;
    #100ns;
  endtask

  task static start_clock();
    fork
      forever begin
        clk_ref_i <= 1;
        #5ns;
        clk_ref_i <= 0;
        #5ns;
      end
    join_none
    @(posedge clk_ref_i);
  endtask

  task static rand_config();
    realtime tick_old;
    realtime tick_new;
    realtime average_timeperiod;
    real fout_exp;
    real fout_got;
    real deviation;
    void'(std::randomize(
        ref_div_i, fb_div_i
    ) with {
      ref_div_i > 0;
      fb_div_i > 0;
      (ref_div_i) <= (100 * fb_div_i);
      (100 * ref_div_i) >= (fb_div_i);
    });
    $display("ref_div_i:%0d\033[20Gfb_div_i:%0d\033[40GFout:%0.3f MHz", ref_div_i, fb_div_i,
             (RefFreq * fb_div_i) / ref_div_i / 1e6);
    do #10ns; while (!locked_o);
    @(posedge clk_o);
    tick_old = $realtime;
    repeat (100) @(posedge clk_o);
    tick_new = $realtime;
    average_timeperiod = (tick_new - tick_old) / 100;
    fout_exp = (RefFreq * fb_div_i) / ref_div_i;
    fout_got = 1s / average_timeperiod;
    deviation = 100 * (fout_got - fout_exp) / fout_exp;
    if (deviation < 0) deviation = -deviation;
    $display("Measured Fout: %0.3f MHz\033[40GTime Period: %0t", 1us / average_timeperiod,
             average_timeperiod);
    $display("Deviation: %0.3f%%\n\n", deviation);


    
    if (deviation > 5) begin
      $display("\033[1;31mERROR: Deviation exceeds 5%%\033[0m");
      test_passed = 0;
    end
  endtask

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-SEQUENTIALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-PROCEDURALS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  initial begin  // main initial

    $dumpfile("pll_tb.vcd");
    $dumpvars(0, pll_tb);
    $timeformat(-9, 2, " ns", 20);

    test_passed = 1;

    apply_reset();
    start_clock();

    repeat (100) rand_config();

    if (test_passed) $display("\033[1;32m************** TEST PASSED **************\033[0m");
    else $display("\033[1;31m************** TEST FAILED **************\033[0m");

    $finish;

  end

endmodule
