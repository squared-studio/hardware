// The decoder_8b10b module is a combinational logic block designed to decode 10-bit input data
// (data_i) into its corresponding 8-bit representation (data_o), adhering to a specific subset of
// the 8b/10b encoding scheme. It also provides a valid_o signal to indicate if the input 10-bit
// code is a recognized valid code.
//
// Author : Foez Ahmed (foez.official@gmail.com)
// This file is part of squared-studio : hardware
// Copyright (c) 2025 squared-studio
// Licensed under the MIT License
// See LICENSE file in the repository root for full license information

module decoder_8b10b (
    input logic [9:0] data_i,  // 10-bit input data to be decoded (8b/10b encoded symbol)

    output logic [7:0] data_o,  // 8-bit decoded output data
    output logic [7:0] k_char_o,  // control character flasg: '1' if data_o is K char, '0' otherwise
    output logic       valid_o    // Output validity flag: '1' if data_i is a valid 8b/10b code, '0' otherwise
);

  //////////////////////////////////////////////////////////////////////////////////////////////////
  //-ASSIGNMENTS
  //////////////////////////////////////////////////////////////////////////////////////////////////

  // Combinational logic to decode the 10-bit input to 8-bit output
  // This 'always_comb' block ensures that outputs update immediately with input changes.
  always_comb begin
    // Case statement to map specific 10-bit 8b/10b encoded patterns to their 8-bit data equivalents.
    // Each line represents a valid 8b/10b code (including both disparities) and its decoded 8-bit value.

    case (data_i)
      10'b1001110100: {data_o, k_char_o, valid_o} = 12'b00000000_0_1;  // D0.0 (RD+)
      10'b0110001011: {data_o, k_char_o, valid_o} = 12'b00000000_0_1;  // D0.0 (RD-)
      10'b0111010100: {data_o, k_char_o, valid_o} = 12'b00000001_0_1;  // D1.0 (RD+)
      10'b1000101011: {data_o, k_char_o, valid_o} = 12'b00000001_0_1;  // D1.0 (RD-)
      10'b1011010100: {data_o, k_char_o, valid_o} = 12'b00000010_0_1;  // D2.0 (RD+)
      10'b0100101011: {data_o, k_char_o, valid_o} = 12'b00000010_0_1;  // D2.0 (RD-)
      10'b1100011011: {data_o, k_char_o, valid_o} = 12'b00000011_0_1;  // D3.0 (RD-)
      10'b1100010100: {data_o, k_char_o, valid_o} = 12'b00000011_0_1;  // D3.0 (RD+)
      10'b1101010100: {data_o, k_char_o, valid_o} = 12'b00000100_0_1;  // D4.0 (RD+)
      10'b0010101011: {data_o, k_char_o, valid_o} = 12'b00000100_0_1;  // D4.0 (RD-)
      10'b1010011011: {data_o, k_char_o, valid_o} = 12'b00000101_0_1;  // D5.0 (RD-)
      10'b1010010100: {data_o, k_char_o, valid_o} = 12'b00000101_0_1;  // D5.0 (RD+)
      10'b0110011011: {data_o, k_char_o, valid_o} = 12'b00000110_0_1;  // D6.0 (RD-)
      10'b0110010100: {data_o, k_char_o, valid_o} = 12'b00000110_0_1;  // D6.0 (RD+)
      10'b1110001011: {data_o, k_char_o, valid_o} = 12'b00000111_0_1;  // D7.0 (RD-)
      10'b0001110100: {data_o, k_char_o, valid_o} = 12'b00000111_0_1;  // D7.0 (RD+)
      10'b1110010100: {data_o, k_char_o, valid_o} = 12'b00001000_0_1;  // D8.0 (RD+)
      10'b0001101011: {data_o, k_char_o, valid_o} = 12'b00001000_0_1;  // D8.0 (RD-)
      10'b1001011011: {data_o, k_char_o, valid_o} = 12'b00001001_0_1;  // D9.0 (RD-)
      10'b1001010100: {data_o, k_char_o, valid_o} = 12'b00001001_0_1;  // D9.0 (RD+)
      10'b0101011011: {data_o, k_char_o, valid_o} = 12'b00001010_0_1;  // D10.0 (RD-)
      10'b0101010100: {data_o, k_char_o, valid_o} = 12'b00001010_0_1;  // D10.0 (RD+)
      10'b1101001011: {data_o, k_char_o, valid_o} = 12'b00001011_0_1;  // D11.0 (RD-)
      10'b1101000100: {data_o, k_char_o, valid_o} = 12'b00001011_0_1;  // D11.0 (RD+)
      10'b0011011011: {data_o, k_char_o, valid_o} = 12'b00001100_0_1;  // D12.0 (RD-)
      10'b0011010100: {data_o, k_char_o, valid_o} = 12'b00001100_0_1;  // D12.0 (RD+)
      10'b1011001011: {data_o, k_char_o, valid_o} = 12'b00001101_0_1;  // D13.0 (RD-)
      10'b1011000100: {data_o, k_char_o, valid_o} = 12'b00001101_0_1;  // D13.0 (RD+)
      10'b0111001011: {data_o, k_char_o, valid_o} = 12'b00001110_0_1;  // D14.0 (RD-)
      10'b0111000100: {data_o, k_char_o, valid_o} = 12'b00001110_0_1;  // D14.0 (RD+)
      10'b0101110100: {data_o, k_char_o, valid_o} = 12'b00001111_0_1;  // D15.0 (RD+)
      10'b1010001011: {data_o, k_char_o, valid_o} = 12'b00001111_0_1;  // D15.0 (RD-)
      10'b0110110100: {data_o, k_char_o, valid_o} = 12'b00010000_0_1;  // D16.0 (RD+)
      10'b1001001011: {data_o, k_char_o, valid_o} = 12'b00010000_0_1;  // D16.0 (RD-)
      10'b1000111011: {data_o, k_char_o, valid_o} = 12'b00010001_0_1;  // D17.0 (RD-)
      10'b1000110100: {data_o, k_char_o, valid_o} = 12'b00010001_0_1;  // D17.0 (RD+)
      10'b0100111011: {data_o, k_char_o, valid_o} = 12'b00010010_0_1;  // D18.0 (RD-)
      10'b0100110100: {data_o, k_char_o, valid_o} = 12'b00010010_0_1;  // D18.0 (RD+)
      10'b1100101011: {data_o, k_char_o, valid_o} = 12'b00010011_0_1;  // D19.0 (RD-)
      10'b1100100100: {data_o, k_char_o, valid_o} = 12'b00010011_0_1;  // D19.0 (RD+)
      10'b0010111011: {data_o, k_char_o, valid_o} = 12'b00010100_0_1;  // D20.0 (RD-)
      10'b0010110100: {data_o, k_char_o, valid_o} = 12'b00010100_0_1;  // D20.0 (RD+)
      10'b1010101011: {data_o, k_char_o, valid_o} = 12'b00010101_0_1;  // D21.0 (RD-)
      10'b1010100100: {data_o, k_char_o, valid_o} = 12'b00010101_0_1;  // D21.0 (RD+)
      10'b0110101011: {data_o, k_char_o, valid_o} = 12'b00010110_0_1;  // D22.0 (RD-)
      10'b0110100100: {data_o, k_char_o, valid_o} = 12'b00010110_0_1;  // D22.0 (RD+)
      10'b1110100100: {data_o, k_char_o, valid_o} = 12'b00010111_0_1;  // D23.0 (RD+)
      10'b0001011011: {data_o, k_char_o, valid_o} = 12'b00010111_0_1;  // D23.0 (RD-)
      10'b1100110100: {data_o, k_char_o, valid_o} = 12'b00011000_0_1;  // D24.0 (RD+)
      10'b0011001011: {data_o, k_char_o, valid_o} = 12'b00011000_0_1;  // D24.0 (RD-)
      10'b1001101011: {data_o, k_char_o, valid_o} = 12'b00011001_0_1;  // D25.0 (RD-)
      10'b1001100100: {data_o, k_char_o, valid_o} = 12'b00011001_0_1;  // D25.0 (RD+)
      10'b0101101011: {data_o, k_char_o, valid_o} = 12'b00011010_0_1;  // D26.0 (RD-)
      10'b0101100100: {data_o, k_char_o, valid_o} = 12'b00011010_0_1;  // D26.0 (RD+)
      10'b1101100100: {data_o, k_char_o, valid_o} = 12'b00011011_0_1;  // D27.0 (RD+)
      10'b0010011011: {data_o, k_char_o, valid_o} = 12'b00011011_0_1;  // D27.0 (RD-)
      10'b0011101011: {data_o, k_char_o, valid_o} = 12'b00011100_0_1;  // D28.0 (RD-)
      10'b0011100100: {data_o, k_char_o, valid_o} = 12'b00011100_0_1;  // D28.0 (RD+)
      10'b1011100100: {data_o, k_char_o, valid_o} = 12'b00011101_0_1;  // D29.0 (RD+)
      10'b0100011011: {data_o, k_char_o, valid_o} = 12'b00011101_0_1;  // D29.0 (RD-)
      10'b0111100100: {data_o, k_char_o, valid_o} = 12'b00011110_0_1;  // D30.0 (RD+)
      10'b1000011011: {data_o, k_char_o, valid_o} = 12'b00011110_0_1;  // D30.0 (RD-)
      10'b1010110100: {data_o, k_char_o, valid_o} = 12'b00011111_0_1;  // D31.0 (RD+)
      10'b0101001011: {data_o, k_char_o, valid_o} = 12'b00011111_0_1;  // D31.0 (RD-)
      10'b1001111001: {data_o, k_char_o, valid_o} = 12'b00100000_0_1;  // D0.1 (RD+)
      10'b0110001001: {data_o, k_char_o, valid_o} = 12'b00100000_0_1;  // D0.1 (RD-)
      10'b0111011001: {data_o, k_char_o, valid_o} = 12'b00100001_0_1;  // D1.1 (RD+)
      10'b1000101001: {data_o, k_char_o, valid_o} = 12'b00100001_0_1;  // D1.1 (RD-)
      10'b1011011001: {data_o, k_char_o, valid_o} = 12'b00100010_0_1;  // D2.1 (RD+)
      10'b0100101001: {data_o, k_char_o, valid_o} = 12'b00100010_0_1;  // D2.1 (RD-)
      10'b1100011001: {data_o, k_char_o, valid_o} = 12'b00100011_0_1;  // D3.1 (RD-)
      10'b1101011001: {data_o, k_char_o, valid_o} = 12'b00100100_0_1;  // D4.1 (RD+)
      10'b0010101001: {data_o, k_char_o, valid_o} = 12'b00100100_0_1;  // D4.1 (RD-)
      10'b1010011001: {data_o, k_char_o, valid_o} = 12'b00100101_0_1;  // D5.1 (RD-)
      10'b0110011001: {data_o, k_char_o, valid_o} = 12'b00100110_0_1;  // D6.1 (RD-)
      10'b1110001001: {data_o, k_char_o, valid_o} = 12'b00100111_0_1;  // D7.1 (RD-)
      10'b0001111001: {data_o, k_char_o, valid_o} = 12'b00100111_0_1;  // D7.1 (RD+)
      10'b1110011001: {data_o, k_char_o, valid_o} = 12'b00101000_0_1;  // D8.1 (RD+)
      10'b0001101001: {data_o, k_char_o, valid_o} = 12'b00101000_0_1;  // D8.1 (RD-)
      10'b1001011001: {data_o, k_char_o, valid_o} = 12'b00101001_0_1;  // D9.1 (RD-)
      10'b0101011001: {data_o, k_char_o, valid_o} = 12'b00101010_0_1;  // D10.1 (RD-)
      10'b1101001001: {data_o, k_char_o, valid_o} = 12'b00101011_0_1;  // D11.1 (RD-)
      10'b0011011001: {data_o, k_char_o, valid_o} = 12'b00101100_0_1;  // D12.1 (RD-)
      10'b1011001001: {data_o, k_char_o, valid_o} = 12'b00101101_0_1;  // D13.1 (RD-)
      10'b0111001001: {data_o, k_char_o, valid_o} = 12'b00101110_0_1;  // D14.1 (RD-)
      10'b0101111001: {data_o, k_char_o, valid_o} = 12'b00101111_0_1;  // D15.1 (RD+)
      10'b1010001001: {data_o, k_char_o, valid_o} = 12'b00101111_0_1;  // D15.1 (RD-)
      10'b0110111001: {data_o, k_char_o, valid_o} = 12'b00110000_0_1;  // D16.1 (RD+)
      10'b1001001001: {data_o, k_char_o, valid_o} = 12'b00110000_0_1;  // D16.1 (RD-)
      10'b1000111001: {data_o, k_char_o, valid_o} = 12'b00110001_0_1;  // D17.1 (RD-)
      10'b0100111001: {data_o, k_char_o, valid_o} = 12'b00110010_0_1;  // D18.1 (RD-)
      10'b1100101001: {data_o, k_char_o, valid_o} = 12'b00110011_0_1;  // D19.1 (RD-)
      10'b0010111001: {data_o, k_char_o, valid_o} = 12'b00110100_0_1;  // D20.1 (RD-)
      10'b1010101001: {data_o, k_char_o, valid_o} = 12'b00110101_0_1;  // D21.1 (RD-)
      10'b0110101001: {data_o, k_char_o, valid_o} = 12'b00110110_0_1;  // D22.1 (RD-)
      10'b1110101001: {data_o, k_char_o, valid_o} = 12'b00110111_0_1;  // D23.1 (RD+)
      10'b0001011001: {data_o, k_char_o, valid_o} = 12'b00110111_0_1;  // D23.1 (RD-)
      10'b1100111001: {data_o, k_char_o, valid_o} = 12'b00111000_0_1;  // D24.1 (RD+)
      10'b0011001001: {data_o, k_char_o, valid_o} = 12'b00111000_0_1;  // D24.1 (RD-)
      10'b1001101001: {data_o, k_char_o, valid_o} = 12'b00111001_0_1;  // D25.1 (RD-)
      10'b0101101001: {data_o, k_char_o, valid_o} = 12'b00111010_0_1;  // D26.1 (RD-)
      10'b1101101001: {data_o, k_char_o, valid_o} = 12'b00111011_0_1;  // D27.1 (RD+)
      10'b0010011001: {data_o, k_char_o, valid_o} = 12'b00111011_0_1;  // D27.1 (RD-)
      10'b0011101001: {data_o, k_char_o, valid_o} = 12'b00111100_0_1;  // D28.1 (RD-)
      10'b1011101001: {data_o, k_char_o, valid_o} = 12'b00111101_0_1;  // D29.1 (RD+)
      10'b0100011001: {data_o, k_char_o, valid_o} = 12'b00111101_0_1;  // D29.1 (RD-)
      10'b0111101001: {data_o, k_char_o, valid_o} = 12'b00111110_0_1;  // D30.1 (RD+)
      10'b1000011001: {data_o, k_char_o, valid_o} = 12'b00111110_0_1;  // D30.1 (RD-)
      10'b1010111001: {data_o, k_char_o, valid_o} = 12'b00111111_0_1;  // D31.1 (RD+)
      10'b0101001001: {data_o, k_char_o, valid_o} = 12'b00111111_0_1;  // D31.1 (RD-)
      10'b1001110101: {data_o, k_char_o, valid_o} = 12'b01000000_0_1;  // D0.2 (RD+)
      10'b0110000101: {data_o, k_char_o, valid_o} = 12'b01000000_0_1;  // D0.2 (RD-)
      10'b0111010101: {data_o, k_char_o, valid_o} = 12'b01000001_0_1;  // D1.2 (RD+)
      10'b1000100101: {data_o, k_char_o, valid_o} = 12'b01000001_0_1;  // D1.2 (RD-)
      10'b1011010101: {data_o, k_char_o, valid_o} = 12'b01000010_0_1;  // D2.2 (RD+)
      10'b0100100101: {data_o, k_char_o, valid_o} = 12'b01000010_0_1;  // D2.2 (RD-)
      10'b1100010101: {data_o, k_char_o, valid_o} = 12'b01000011_0_1;  // D3.2 (RD+)
      10'b1101010101: {data_o, k_char_o, valid_o} = 12'b01000100_0_1;  // D4.2 (RD+)
      10'b0010100101: {data_o, k_char_o, valid_o} = 12'b01000100_0_1;  // D4.2 (RD-)
      10'b1010010101: {data_o, k_char_o, valid_o} = 12'b01000101_0_1;  // D5.2 (RD+)
      10'b0110010101: {data_o, k_char_o, valid_o} = 12'b01000110_0_1;  // D6.2 (RD+)
      10'b1110000101: {data_o, k_char_o, valid_o} = 12'b01000111_0_1;  // D7.2 (RD+)
      10'b0001110101: {data_o, k_char_o, valid_o} = 12'b01000111_0_1;  // D7.2 (RD-)
      10'b1110010101: {data_o, k_char_o, valid_o} = 12'b01001000_0_1;  // D8.2 (RD+)
      10'b0001100101: {data_o, k_char_o, valid_o} = 12'b01001000_0_1;  // D8.2 (RD-)
      10'b1001010101: {data_o, k_char_o, valid_o} = 12'b01001001_0_1;  // D9.2 (RD+)
      10'b0101010101: {data_o, k_char_o, valid_o} = 12'b01001010_0_1;  // D10.2 (RD+)
      10'b1101000101: {data_o, k_char_o, valid_o} = 12'b01001011_0_1;  // D11.2 (RD+)
      10'b0011010101: {data_o, k_char_o, valid_o} = 12'b01001100_0_1;  // D12.2 (RD+)
      10'b1011000101: {data_o, k_char_o, valid_o} = 12'b01001101_0_1;  // D13.2 (RD+)
      10'b0111000101: {data_o, k_char_o, valid_o} = 12'b01001110_0_1;  // D14.2 (RD+)
      10'b0101110101: {data_o, k_char_o, valid_o} = 12'b01001111_0_1;  // D15.2 (RD+)
      10'b1010000101: {data_o, k_char_o, valid_o} = 12'b01001111_0_1;  // D15.2 (RD-)
      10'b0110110101: {data_o, k_char_o, valid_o} = 12'b01010000_0_1;  // D16.2 (RD+)
      10'b1001000101: {data_o, k_char_o, valid_o} = 12'b01010000_0_1;  // D16.2 (RD-)
      10'b1000110101: {data_o, k_char_o, valid_o} = 12'b01010001_0_1;  // D17.2 (RD+)
      10'b0100110101: {data_o, k_char_o, valid_o} = 12'b01010010_0_1;  // D18.2 (RD+)
      10'b1100100101: {data_o, k_char_o, valid_o} = 12'b01010011_0_1;  // D19.2 (RD+)
      10'b0010110101: {data_o, k_char_o, valid_o} = 12'b01010100_0_1;  // D20.2 (RD+)
      10'b1010100101: {data_o, k_char_o, valid_o} = 12'b01010101_0_1;  // D21.2 (RD+)
      10'b0110100101: {data_o, k_char_o, valid_o} = 12'b01010110_0_1;  // D22.2 (RD+)
      10'b1110100101: {data_o, k_char_o, valid_o} = 12'b01010111_0_1;  // D23.2 (RD+)
      10'b0001010101: {data_o, k_char_o, valid_o} = 12'b01010111_0_1;  // D23.2 (RD-)
      10'b1100110101: {data_o, k_char_o, valid_o} = 12'b01011000_0_1;  // D24.2 (RD+)
      10'b0011000101: {data_o, k_char_o, valid_o} = 12'b01011000_0_1;  // D24.2 (RD-)
      10'b1001100101: {data_o, k_char_o, valid_o} = 12'b01011001_0_1;  // D25.2 (RD+)
      10'b0101100101: {data_o, k_char_o, valid_o} = 12'b01011010_0_1;  // D26.2 (RD+)
      10'b1101100101: {data_o, k_char_o, valid_o} = 12'b01011011_0_1;  // D27.2 (RD+)
      10'b0010010101: {data_o, k_char_o, valid_o} = 12'b01011011_0_1;  // D27.2 (RD-)
      10'b0011100101: {data_o, k_char_o, valid_o} = 12'b01011100_0_1;  // D28.2 (RD+)
      10'b1011100101: {data_o, k_char_o, valid_o} = 12'b01011101_0_1;  // D29.2 (RD+)
      10'b0100010101: {data_o, k_char_o, valid_o} = 12'b01011101_0_1;  // D29.2 (RD-)
      10'b0111100101: {data_o, k_char_o, valid_o} = 12'b01011110_0_1;  // D30.2 (RD+)
      10'b1000010101: {data_o, k_char_o, valid_o} = 12'b01011110_0_1;  // D30.2 (RD-)
      10'b1010110101: {data_o, k_char_o, valid_o} = 12'b01011111_0_1;  // D31.2 (RD+)
      10'b0101000101: {data_o, k_char_o, valid_o} = 12'b01011111_0_1;  // D31.2 (RD-)
      10'b1001110011: {data_o, k_char_o, valid_o} = 12'b01100000_0_1;  // D0.3 (RD+)
      10'b0110001100: {data_o, k_char_o, valid_o} = 12'b01100000_0_1;  // D0.3 (RD-)
      10'b0111010011: {data_o, k_char_o, valid_o} = 12'b01100001_0_1;  // D1.3 (RD+)
      10'b1000101100: {data_o, k_char_o, valid_o} = 12'b01100001_0_1;  // D1.3 (RD-)
      10'b1011010011: {data_o, k_char_o, valid_o} = 12'b01100010_0_1;  // D2.3 (RD+)
      10'b0100101100: {data_o, k_char_o, valid_o} = 12'b01100010_0_1;  // D2.3 (RD-)
      10'b1100011100: {data_o, k_char_o, valid_o} = 12'b01100011_0_1;  // D3.3 (RD-)
      10'b1100010011: {data_o, k_char_o, valid_o} = 12'b01100011_0_1;  // D3.3 (RD+)
      10'b1101010011: {data_o, k_char_o, valid_o} = 12'b01100100_0_1;  // D4.3 (RD+)
      10'b0010101100: {data_o, k_char_o, valid_o} = 12'b01100100_0_1;  // D4.3 (RD-)
      10'b1010011100: {data_o, k_char_o, valid_o} = 12'b01100101_0_1;  // D5.3 (RD-)
      10'b1010010011: {data_o, k_char_o, valid_o} = 12'b01100101_0_1;  // D5.3 (RD+)
      10'b0110011100: {data_o, k_char_o, valid_o} = 12'b01100110_0_1;  // D6.3 (RD-)
      10'b0110010011: {data_o, k_char_o, valid_o} = 12'b01100110_0_1;  // D6.3 (RD+)
      10'b1110001100: {data_o, k_char_o, valid_o} = 12'b01100111_0_1;  // D7.3 (RD-)
      10'b0001110011: {data_o, k_char_o, valid_o} = 12'b01100111_0_1;  // D7.3 (RD+)
      10'b1110010011: {data_o, k_char_o, valid_o} = 12'b01101000_0_1;  // D8.3 (RD+)
      10'b0001101100: {data_o, k_char_o, valid_o} = 12'b01101000_0_1;  // D8.3 (RD-)
      10'b1001011100: {data_o, k_char_o, valid_o} = 12'b01101001_0_1;  // D9.3 (RD-)
      10'b1001010011: {data_o, k_char_o, valid_o} = 12'b01101001_0_1;  // D9.3 (RD+)
      10'b0101011100: {data_o, k_char_o, valid_o} = 12'b01101010_0_1;  // D10.3 (RD-)
      10'b0101010011: {data_o, k_char_o, valid_o} = 12'b01101010_0_1;  // D10.3 (RD+)
      10'b1101001100: {data_o, k_char_o, valid_o} = 12'b01101011_0_1;  // D11.3 (RD-)
      10'b1101000011: {data_o, k_char_o, valid_o} = 12'b01101011_0_1;  // D11.3 (RD+)
      10'b0011011100: {data_o, k_char_o, valid_o} = 12'b01101100_0_1;  // D12.3 (RD-)
      10'b0011010011: {data_o, k_char_o, valid_o} = 12'b01101100_0_1;  // D12.3 (RD+)
      10'b1011001100: {data_o, k_char_o, valid_o} = 12'b01101101_0_1;  // D13.3 (RD-)
      10'b1011000011: {data_o, k_char_o, valid_o} = 12'b01101101_0_1;  // D13.3 (RD+)
      10'b0111001100: {data_o, k_char_o, valid_o} = 12'b01101110_0_1;  // D14.3 (RD-)
      10'b0111000011: {data_o, k_char_o, valid_o} = 12'b01101110_0_1;  // D14.3 (RD+)
      10'b0101110011: {data_o, k_char_o, valid_o} = 12'b01101111_0_1;  // D15.3 (RD+)
      10'b1010001100: {data_o, k_char_o, valid_o} = 12'b01101111_0_1;  // D15.3 (RD-)
      10'b0110110011: {data_o, k_char_o, valid_o} = 12'b01110000_0_1;  // D16.3 (RD+)
      10'b1001001100: {data_o, k_char_o, valid_o} = 12'b01110000_0_1;  // D16.3 (RD-)
      10'b1000111100: {data_o, k_char_o, valid_o} = 12'b01110001_0_1;  // D17.3 (RD-)
      10'b1000110011: {data_o, k_char_o, valid_o} = 12'b01110001_0_1;  // D17.3 (RD+)
      10'b0100111100: {data_o, k_char_o, valid_o} = 12'b01110010_0_1;  // D18.3 (RD-)
      10'b0100110011: {data_o, k_char_o, valid_o} = 12'b01110010_0_1;  // D18.3 (RD+)
      10'b1100101100: {data_o, k_char_o, valid_o} = 12'b01110011_0_1;  // D19.3 (RD-)
      10'b1100100011: {data_o, k_char_o, valid_o} = 12'b01110011_0_1;  // D19.3 (RD+)
      10'b0010111100: {data_o, k_char_o, valid_o} = 12'b01110100_0_1;  // D20.3 (RD-)
      10'b0010110011: {data_o, k_char_o, valid_o} = 12'b01110100_0_1;  // D20.3 (RD+)
      10'b1010101100: {data_o, k_char_o, valid_o} = 12'b01110101_0_1;  // D21.3 (RD-)
      10'b1010100011: {data_o, k_char_o, valid_o} = 12'b01110101_0_1;  // D21.3 (RD+)
      10'b0110101100: {data_o, k_char_o, valid_o} = 12'b01110110_0_1;  // D22.3 (RD-)
      10'b0110100011: {data_o, k_char_o, valid_o} = 12'b01110110_0_1;  // D22.3 (RD+)
      10'b1110100011: {data_o, k_char_o, valid_o} = 12'b01110111_0_1;  // D23.3 (RD+)
      10'b0001011100: {data_o, k_char_o, valid_o} = 12'b01110111_0_1;  // D23.3 (RD-)
      10'b1100110011: {data_o, k_char_o, valid_o} = 12'b01111000_0_1;  // D24.3 (RD+)
      10'b0011001100: {data_o, k_char_o, valid_o} = 12'b01111000_0_1;  // D24.3 (RD-)
      10'b1001101100: {data_o, k_char_o, valid_o} = 12'b01111001_0_1;  // D25.3 (RD-)
      10'b1001100011: {data_o, k_char_o, valid_o} = 12'b01111001_0_1;  // D25.3 (RD+)
      10'b0101101100: {data_o, k_char_o, valid_o} = 12'b01111010_0_1;  // D26.3 (RD-)
      10'b0101100011: {data_o, k_char_o, valid_o} = 12'b01111010_0_1;  // D26.3 (RD+)
      10'b1101100011: {data_o, k_char_o, valid_o} = 12'b01111011_0_1;  // D27.3 (RD+)
      10'b0010011100: {data_o, k_char_o, valid_o} = 12'b01111011_0_1;  // D27.3 (RD-)
      10'b0011101100: {data_o, k_char_o, valid_o} = 12'b01111100_0_1;  // D28.3 (RD-)
      10'b0011100011: {data_o, k_char_o, valid_o} = 12'b01111100_0_1;  // D28.3 (RD+)
      10'b1011100011: {data_o, k_char_o, valid_o} = 12'b01111101_0_1;  // D29.3 (RD+)
      10'b0100011100: {data_o, k_char_o, valid_o} = 12'b01111101_0_1;  // D29.3 (RD-)
      10'b0111100011: {data_o, k_char_o, valid_o} = 12'b01111110_0_1;  // D30.3 (RD+)
      10'b1000011100: {data_o, k_char_o, valid_o} = 12'b01111110_0_1;  // D30.3 (RD-)
      10'b1010110011: {data_o, k_char_o, valid_o} = 12'b01111111_0_1;  // D31.3 (RD+)
      10'b0101001100: {data_o, k_char_o, valid_o} = 12'b01111111_0_1;  // D31.3 (RD-)
      10'b1001110010: {data_o, k_char_o, valid_o} = 12'b10000000_0_1;  // D0.4 (RD+)
      10'b0110001101: {data_o, k_char_o, valid_o} = 12'b10000000_0_1;  // D0.4 (RD-)
      10'b0111010010: {data_o, k_char_o, valid_o} = 12'b10000001_0_1;  // D1.4 (RD+)
      10'b1000101101: {data_o, k_char_o, valid_o} = 12'b10000001_0_1;  // D1.4 (RD-)
      10'b1011010010: {data_o, k_char_o, valid_o} = 12'b10000010_0_1;  // D2.4 (RD+)
      10'b0100101101: {data_o, k_char_o, valid_o} = 12'b10000010_0_1;  // D2.4 (RD-)
      10'b1100011101: {data_o, k_char_o, valid_o} = 12'b10000011_0_1;  // D3.4 (RD-)
      10'b1100010010: {data_o, k_char_o, valid_o} = 12'b10000011_0_1;  // D3.4 (RD+)
      10'b1101010010: {data_o, k_char_o, valid_o} = 12'b10000100_0_1;  // D4.4 (RD+)
      10'b0010101101: {data_o, k_char_o, valid_o} = 12'b10000100_0_1;  // D4.4 (RD-)
      10'b1010011101: {data_o, k_char_o, valid_o} = 12'b10000101_0_1;  // D5.4 (RD-)
      10'b1010010010: {data_o, k_char_o, valid_o} = 12'b10000101_0_1;  // D5.4 (RD+)
      10'b0110011101: {data_o, k_char_o, valid_o} = 12'b10000110_0_1;  // D6.4 (RD-)
      10'b0110010010: {data_o, k_char_o, valid_o} = 12'b10000110_0_1;  // D6.4 (RD+)
      10'b1110001101: {data_o, k_char_o, valid_o} = 12'b10000111_0_1;  // D7.4 (RD-)
      10'b0001110010: {data_o, k_char_o, valid_o} = 12'b10000111_0_1;  // D7.4 (RD+)
      10'b1110010010: {data_o, k_char_o, valid_o} = 12'b10001000_0_1;  // D8.4 (RD+)
      10'b0001101101: {data_o, k_char_o, valid_o} = 12'b10001000_0_1;  // D8.4 (RD-)
      10'b1001011101: {data_o, k_char_o, valid_o} = 12'b10001001_0_1;  // D9.4 (RD-)
      10'b1001010010: {data_o, k_char_o, valid_o} = 12'b10001001_0_1;  // D9.4 (RD+)
      10'b0101011101: {data_o, k_char_o, valid_o} = 12'b10001010_0_1;  // D10.4 (RD-)
      10'b0101010010: {data_o, k_char_o, valid_o} = 12'b10001010_0_1;  // D10.4 (RD+)
      10'b1101001101: {data_o, k_char_o, valid_o} = 12'b10001011_0_1;  // D11.4 (RD-)
      10'b1101000010: {data_o, k_char_o, valid_o} = 12'b10001011_0_1;  // D11.4 (RD+)
      10'b0011011101: {data_o, k_char_o, valid_o} = 12'b10001100_0_1;  // D12.4 (RD-)
      10'b0011010010: {data_o, k_char_o, valid_o} = 12'b10001100_0_1;  // D12.4 (RD+)
      10'b1011001101: {data_o, k_char_o, valid_o} = 12'b10001101_0_1;  // D13.4 (RD-)
      10'b1011000010: {data_o, k_char_o, valid_o} = 12'b10001101_0_1;  // D13.4 (RD+)
      10'b0111001101: {data_o, k_char_o, valid_o} = 12'b10001110_0_1;  // D14.4 (RD-)
      10'b0111000010: {data_o, k_char_o, valid_o} = 12'b10001110_0_1;  // D14.4 (RD+)
      10'b0101110010: {data_o, k_char_o, valid_o} = 12'b10001111_0_1;  // D15.4 (RD+)
      10'b1010001101: {data_o, k_char_o, valid_o} = 12'b10001111_0_1;  // D15.4 (RD-)
      10'b0110110010: {data_o, k_char_o, valid_o} = 12'b10010000_0_1;  // D16.4 (RD+)
      10'b1001001101: {data_o, k_char_o, valid_o} = 12'b10010000_0_1;  // D16.4 (RD-)
      10'b1000111101: {data_o, k_char_o, valid_o} = 12'b10010001_0_1;  // D17.4 (RD-)
      10'b1000110010: {data_o, k_char_o, valid_o} = 12'b10010001_0_1;  // D17.4 (RD+)
      10'b0100111101: {data_o, k_char_o, valid_o} = 12'b10010010_0_1;  // D18.4 (RD-)
      10'b0100110010: {data_o, k_char_o, valid_o} = 12'b10010010_0_1;  // D18.4 (RD+)
      10'b1100101101: {data_o, k_char_o, valid_o} = 12'b10010011_0_1;  // D19.4 (RD-)
      10'b1100100010: {data_o, k_char_o, valid_o} = 12'b10010011_0_1;  // D19.4 (RD+)
      10'b0010111101: {data_o, k_char_o, valid_o} = 12'b10010100_0_1;  // D20.4 (RD-)
      10'b0010110010: {data_o, k_char_o, valid_o} = 12'b10010100_0_1;  // D20.4 (RD+)
      10'b1010101101: {data_o, k_char_o, valid_o} = 12'b10010101_0_1;  // D21.4 (RD-)
      10'b1010100010: {data_o, k_char_o, valid_o} = 12'b10010101_0_1;  // D21.4 (RD+)
      10'b0110101101: {data_o, k_char_o, valid_o} = 12'b10010110_0_1;  // D22.4 (RD-)
      10'b0110100010: {data_o, k_char_o, valid_o} = 12'b10010110_0_1;  // D22.4 (RD+)
      10'b1110100010: {data_o, k_char_o, valid_o} = 12'b10010111_0_1;  // D23.4 (RD+)
      10'b0001011101: {data_o, k_char_o, valid_o} = 12'b10010111_0_1;  // D23.4 (RD-)
      10'b1100110010: {data_o, k_char_o, valid_o} = 12'b10011000_0_1;  // D24.4 (RD+)
      10'b0011001101: {data_o, k_char_o, valid_o} = 12'b10011000_0_1;  // D24.4 (RD-)
      10'b1001101101: {data_o, k_char_o, valid_o} = 12'b10011001_0_1;  // D25.4 (RD-)
      10'b1001100010: {data_o, k_char_o, valid_o} = 12'b10011001_0_1;  // D25.4 (RD+)
      10'b0101101101: {data_o, k_char_o, valid_o} = 12'b10011010_0_1;  // D26.4 (RD-)
      10'b0101100010: {data_o, k_char_o, valid_o} = 12'b10011010_0_1;  // D26.4 (RD+)
      10'b1101100010: {data_o, k_char_o, valid_o} = 12'b10011011_0_1;  // D27.4 (RD+)
      10'b0010011101: {data_o, k_char_o, valid_o} = 12'b10011011_0_1;  // D27.4 (RD-)
      10'b0011101101: {data_o, k_char_o, valid_o} = 12'b10011100_0_1;  // D28.4 (RD-)
      10'b0011100010: {data_o, k_char_o, valid_o} = 12'b10011100_0_1;  // D28.4 (RD+)
      10'b1011100010: {data_o, k_char_o, valid_o} = 12'b10011101_0_1;  // D29.4 (RD+)
      10'b0100011101: {data_o, k_char_o, valid_o} = 12'b10011101_0_1;  // D29.4 (RD-)
      10'b0111100010: {data_o, k_char_o, valid_o} = 12'b10011110_0_1;  // D30.4 (RD+)
      10'b1000011101: {data_o, k_char_o, valid_o} = 12'b10011110_0_1;  // D30.4 (RD-)
      10'b1010110010: {data_o, k_char_o, valid_o} = 12'b10011111_0_1;  // D31.4 (RD+)
      10'b0101001101: {data_o, k_char_o, valid_o} = 12'b10011111_0_1;  // D31.4 (RD-)
      10'b1001111010: {data_o, k_char_o, valid_o} = 12'b10100000_0_1;  // D0.5 (RD+)
      10'b0110001010: {data_o, k_char_o, valid_o} = 12'b10100000_0_1;  // D0.5 (RD-)
      10'b0111011010: {data_o, k_char_o, valid_o} = 12'b10100001_0_1;  // D1.5 (RD+)
      10'b1000101010: {data_o, k_char_o, valid_o} = 12'b10100001_0_1;  // D1.5 (RD-)
      10'b1011011010: {data_o, k_char_o, valid_o} = 12'b10100010_0_1;  // D2.5 (RD+)
      10'b0100101010: {data_o, k_char_o, valid_o} = 12'b10100010_0_1;  // D2.5 (RD-)
      10'b1100011010: {data_o, k_char_o, valid_o} = 12'b10100011_0_1;  // D3.5 (RD-)
      10'b1101011010: {data_o, k_char_o, valid_o} = 12'b10100100_0_1;  // D4.5 (RD+)
      10'b0010101010: {data_o, k_char_o, valid_o} = 12'b10100100_0_1;  // D4.5 (RD-)
      10'b1010011010: {data_o, k_char_o, valid_o} = 12'b10100101_0_1;  // D5.5 (RD-)
      10'b0110011010: {data_o, k_char_o, valid_o} = 12'b10100110_0_1;  // D6.5 (RD-)
      10'b1110001010: {data_o, k_char_o, valid_o} = 12'b10100111_0_1;  // D7.5 (RD-)
      10'b0001111010: {data_o, k_char_o, valid_o} = 12'b10100111_0_1;  // D7.5 (RD+)
      10'b1110011010: {data_o, k_char_o, valid_o} = 12'b10101000_0_1;  // D8.5 (RD+)
      10'b0001101010: {data_o, k_char_o, valid_o} = 12'b10101000_0_1;  // D8.5 (RD-)
      10'b1001011010: {data_o, k_char_o, valid_o} = 12'b10101001_0_1;  // D9.5 (RD-)
      10'b0101011010: {data_o, k_char_o, valid_o} = 12'b10101010_0_1;  // D10.5 (RD-)
      10'b1101001010: {data_o, k_char_o, valid_o} = 12'b10101011_0_1;  // D11.5 (RD-)
      10'b0011011010: {data_o, k_char_o, valid_o} = 12'b10101100_0_1;  // D12.5 (RD-)
      10'b1011001010: {data_o, k_char_o, valid_o} = 12'b10101101_0_1;  // D13.5 (RD-)
      10'b0111001010: {data_o, k_char_o, valid_o} = 12'b10101110_0_1;  // D14.5 (RD-)
      10'b0101111010: {data_o, k_char_o, valid_o} = 12'b10101111_0_1;  // D15.5 (RD+)
      10'b1010001010: {data_o, k_char_o, valid_o} = 12'b10101111_0_1;  // D15.5 (RD-)
      10'b0110111010: {data_o, k_char_o, valid_o} = 12'b10110000_0_1;  // D16.5 (RD+)
      10'b1001001010: {data_o, k_char_o, valid_o} = 12'b10110000_0_1;  // D16.5 (RD-)
      10'b1000111010: {data_o, k_char_o, valid_o} = 12'b10110001_0_1;  // D17.5 (RD-)
      10'b0100111010: {data_o, k_char_o, valid_o} = 12'b10110010_0_1;  // D18.5 (RD-)
      10'b1100101010: {data_o, k_char_o, valid_o} = 12'b10110011_0_1;  // D19.5 (RD-)
      10'b0010111010: {data_o, k_char_o, valid_o} = 12'b10110100_0_1;  // D20.5 (RD-)
      10'b1010101010: {data_o, k_char_o, valid_o} = 12'b10110101_0_1;  // D21.5 (RD-)
      10'b0110101010: {data_o, k_char_o, valid_o} = 12'b10110110_0_1;  // D22.5 (RD-)
      10'b1110101010: {data_o, k_char_o, valid_o} = 12'b10110111_0_1;  // D23.5 (RD+)
      10'b0001011010: {data_o, k_char_o, valid_o} = 12'b10110111_0_1;  // D23.5 (RD-)
      10'b1100111010: {data_o, k_char_o, valid_o} = 12'b10111000_0_1;  // D24.5 (RD+)
      10'b0011001010: {data_o, k_char_o, valid_o} = 12'b10111000_0_1;  // D24.5 (RD-)
      10'b1001101010: {data_o, k_char_o, valid_o} = 12'b10111001_0_1;  // D25.5 (RD-)
      10'b0101101010: {data_o, k_char_o, valid_o} = 12'b10111010_0_1;  // D26.5 (RD-)
      10'b1101101010: {data_o, k_char_o, valid_o} = 12'b10111011_0_1;  // D27.5 (RD+)
      10'b0010011010: {data_o, k_char_o, valid_o} = 12'b10111011_0_1;  // D27.5 (RD-)
      10'b0011101010: {data_o, k_char_o, valid_o} = 12'b10111100_0_1;  // D28.5 (RD-)
      10'b1011101010: {data_o, k_char_o, valid_o} = 12'b10111101_0_1;  // D29.5 (RD+)
      10'b0100011010: {data_o, k_char_o, valid_o} = 12'b10111101_0_1;  // D29.5 (RD-)
      10'b0111101010: {data_o, k_char_o, valid_o} = 12'b10111110_0_1;  // D30.5 (RD+)
      10'b1000011010: {data_o, k_char_o, valid_o} = 12'b10111110_0_1;  // D30.5 (RD-)
      10'b1010111010: {data_o, k_char_o, valid_o} = 12'b10111111_0_1;  // D31.5 (RD+)
      10'b0101001010: {data_o, k_char_o, valid_o} = 12'b10111111_0_1;  // D31.5 (RD-)
      10'b1001110110: {data_o, k_char_o, valid_o} = 12'b11000000_0_1;  // D0.6 (RD+)
      10'b0110000110: {data_o, k_char_o, valid_o} = 12'b11000000_0_1;  // D0.6 (RD-)
      10'b0111010110: {data_o, k_char_o, valid_o} = 12'b11000001_0_1;  // D1.6 (RD+)
      10'b1000100110: {data_o, k_char_o, valid_o} = 12'b11000001_0_1;  // D1.6 (RD-)
      10'b1011010110: {data_o, k_char_o, valid_o} = 12'b11000010_0_1;  // D2.6 (RD+)
      10'b0100100110: {data_o, k_char_o, valid_o} = 12'b11000010_0_1;  // D2.6 (RD-)
      10'b1100010110: {data_o, k_char_o, valid_o} = 12'b11000011_0_1;  // D3.6 (RD+)
      10'b1101010110: {data_o, k_char_o, valid_o} = 12'b11000100_0_1;  // D4.6 (RD+)
      10'b0010100110: {data_o, k_char_o, valid_o} = 12'b11000100_0_1;  // D4.6 (RD-)
      10'b1010010110: {data_o, k_char_o, valid_o} = 12'b11000101_0_1;  // D5.6 (RD+)
      10'b0110010110: {data_o, k_char_o, valid_o} = 12'b11000110_0_1;  // D6.6 (RD+)
      10'b1110000110: {data_o, k_char_o, valid_o} = 12'b11000111_0_1;  // D7.6 (RD+)
      10'b0001110110: {data_o, k_char_o, valid_o} = 12'b11000111_0_1;  // D7.6 (RD-)
      10'b1110010110: {data_o, k_char_o, valid_o} = 12'b11001000_0_1;  // D8.6 (RD+)
      10'b0001100110: {data_o, k_char_o, valid_o} = 12'b11001000_0_1;  // D8.6 (RD-)
      10'b1001010110: {data_o, k_char_o, valid_o} = 12'b11001001_0_1;  // D9.6 (RD+)
      10'b0101010110: {data_o, k_char_o, valid_o} = 12'b11001010_0_1;  // D10.6 (RD+)
      10'b1101000110: {data_o, k_char_o, valid_o} = 12'b11001011_0_1;  // D11.6 (RD+)
      10'b0011010110: {data_o, k_char_o, valid_o} = 12'b11001100_0_1;  // D12.6 (RD+)
      10'b1011000110: {data_o, k_char_o, valid_o} = 12'b11001101_0_1;  // D13.6 (RD+)
      10'b0111000110: {data_o, k_char_o, valid_o} = 12'b11001110_0_1;  // D14.6 (RD+)
      10'b0101110110: {data_o, k_char_o, valid_o} = 12'b11001111_0_1;  // D15.6 (RD+)
      10'b1010000110: {data_o, k_char_o, valid_o} = 12'b11001111_0_1;  // D15.6 (RD-)
      10'b0110110110: {data_o, k_char_o, valid_o} = 12'b11010000_0_1;  // D16.6 (RD+)
      10'b1001000110: {data_o, k_char_o, valid_o} = 12'b11010000_0_1;  // D16.6 (RD-)
      10'b1000110110: {data_o, k_char_o, valid_o} = 12'b11010001_0_1;  // D17.6 (RD+)
      10'b0100110110: {data_o, k_char_o, valid_o} = 12'b11010010_0_1;  // D18.6 (RD+)
      10'b1100100110: {data_o, k_char_o, valid_o} = 12'b11010011_0_1;  // D19.6 (RD+)
      10'b0010110110: {data_o, k_char_o, valid_o} = 12'b11010100_0_1;  // D20.6 (RD+)
      10'b1010100110: {data_o, k_char_o, valid_o} = 12'b11010101_0_1;  // D21.6 (RD+)
      10'b0110100110: {data_o, k_char_o, valid_o} = 12'b11010110_0_1;  // D22.6 (RD+)
      10'b1110100110: {data_o, k_char_o, valid_o} = 12'b11010111_0_1;  // D23.6 (RD+)
      10'b0001010110: {data_o, k_char_o, valid_o} = 12'b11010111_0_1;  // D23.6 (RD-)
      10'b1100110110: {data_o, k_char_o, valid_o} = 12'b11011000_0_1;  // D24.6 (RD+)
      10'b0011000110: {data_o, k_char_o, valid_o} = 12'b11011000_0_1;  // D24.6 (RD-)
      10'b1001100110: {data_o, k_char_o, valid_o} = 12'b11011001_0_1;  // D25.6 (RD+)
      10'b0101100110: {data_o, k_char_o, valid_o} = 12'b11011010_0_1;  // D26.6 (RD+)
      10'b1101100110: {data_o, k_char_o, valid_o} = 12'b11011011_0_1;  // D27.6 (RD+)
      10'b0010010110: {data_o, k_char_o, valid_o} = 12'b11011011_0_1;  // D27.6 (RD-)
      10'b0011100110: {data_o, k_char_o, valid_o} = 12'b11011100_0_1;  // D28.6 (RD+)
      10'b1011100110: {data_o, k_char_o, valid_o} = 12'b11011101_0_1;  // D29.6 (RD+)
      10'b0100010110: {data_o, k_char_o, valid_o} = 12'b11011101_0_1;  // D29.6 (RD-)
      10'b0111100110: {data_o, k_char_o, valid_o} = 12'b11011110_0_1;  // D30.6 (RD+)
      10'b1000010110: {data_o, k_char_o, valid_o} = 12'b11011110_0_1;  // D30.6 (RD-)
      10'b1010110110: {data_o, k_char_o, valid_o} = 12'b11011111_0_1;  // D31.6 (RD+)
      10'b0101000110: {data_o, k_char_o, valid_o} = 12'b11011111_0_1;  // D31.6 (RD-)
      10'b1001110001: {data_o, k_char_o, valid_o} = 12'b11100000_0_1;  // D0.7 (RD+)
      10'b0110001110: {data_o, k_char_o, valid_o} = 12'b11100000_0_1;  // D0.7 (RD-)
      10'b0111010001: {data_o, k_char_o, valid_o} = 12'b11100001_0_1;  // D1.7 (RD+)
      10'b1000101110: {data_o, k_char_o, valid_o} = 12'b11100001_0_1;  // D1.7 (RD-)
      10'b1011010001: {data_o, k_char_o, valid_o} = 12'b11100010_0_1;  // D2.7 (RD+)
      10'b0100101110: {data_o, k_char_o, valid_o} = 12'b11100010_0_1;  // D2.7 (RD-)
      10'b1100011110: {data_o, k_char_o, valid_o} = 12'b11100011_0_1;  // D3.7 (RD-)
      10'b1100010001: {data_o, k_char_o, valid_o} = 12'b11100011_0_1;  // D3.7 (RD+)
      10'b1101010001: {data_o, k_char_o, valid_o} = 12'b11100100_0_1;  // D4.7 (RD+)
      10'b0010101110: {data_o, k_char_o, valid_o} = 12'b11100100_0_1;  // D4.7 (RD-)
      10'b1010011110: {data_o, k_char_o, valid_o} = 12'b11100101_0_1;  // D5.7 (RD-)
      10'b1010010001: {data_o, k_char_o, valid_o} = 12'b11100101_0_1;  // D5.7 (RD+)
      10'b0110011110: {data_o, k_char_o, valid_o} = 12'b11100110_0_1;  // D6.7 (RD-)
      10'b0110010001: {data_o, k_char_o, valid_o} = 12'b11100110_0_1;  // D6.7 (RD+)
      10'b1110001110: {data_o, k_char_o, valid_o} = 12'b11100111_0_1;  // D7.7 (RD-)
      10'b0001110001: {data_o, k_char_o, valid_o} = 12'b11100111_0_1;  // D7.7 (RD+)
      10'b1110010001: {data_o, k_char_o, valid_o} = 12'b11101000_0_1;  // D8.7 (RD+)
      10'b0001101110: {data_o, k_char_o, valid_o} = 12'b11101000_0_1;  // D8.7 (RD-)
      10'b1001011110: {data_o, k_char_o, valid_o} = 12'b11101001_0_1;  // D9.7 (RD-)
      10'b1001010001: {data_o, k_char_o, valid_o} = 12'b11101001_0_1;  // D9.7 (RD+)
      10'b0101011110: {data_o, k_char_o, valid_o} = 12'b11101010_0_1;  // D10.7 (RD-)
      10'b0101010001: {data_o, k_char_o, valid_o} = 12'b11101010_0_1;  // D10.7 (RD+)
      10'b1101001110: {data_o, k_char_o, valid_o} = 12'b11101011_0_1;  // D11.7 (RD-)
      10'b1101001000: {data_o, k_char_o, valid_o} = 12'b11101011_0_1;  // D11.7 (RD+)
      10'b0011011110: {data_o, k_char_o, valid_o} = 12'b11101100_0_1;  // D12.7 (RD-)
      10'b0011010001: {data_o, k_char_o, valid_o} = 12'b11101100_0_1;  // D12.7 (RD+)
      10'b1011001110: {data_o, k_char_o, valid_o} = 12'b11101101_0_1;  // D13.7 (RD-)
      10'b1011001000: {data_o, k_char_o, valid_o} = 12'b11101101_0_1;  // D13.7 (RD+)
      10'b0111001110: {data_o, k_char_o, valid_o} = 12'b11101110_0_1;  // D14.7 (RD-)
      10'b0111001000: {data_o, k_char_o, valid_o} = 12'b11101110_0_1;  // D14.7 (RD+)
      10'b0101110001: {data_o, k_char_o, valid_o} = 12'b11101111_0_1;  // D15.7 (RD+)
      10'b1010001110: {data_o, k_char_o, valid_o} = 12'b11101111_0_1;  // D15.7 (RD-)
      10'b0110110001: {data_o, k_char_o, valid_o} = 12'b11110000_0_1;  // D16.7 (RD+)
      10'b1001001110: {data_o, k_char_o, valid_o} = 12'b11110000_0_1;  // D16.7 (RD-)
      10'b1000110111: {data_o, k_char_o, valid_o} = 12'b11110001_0_1;  // D17.7 (RD-)
      10'b1000110001: {data_o, k_char_o, valid_o} = 12'b11110001_0_1;  // D17.7 (RD+)
      10'b0100110111: {data_o, k_char_o, valid_o} = 12'b11110010_0_1;  // D18.7 (RD-)
      10'b0100110001: {data_o, k_char_o, valid_o} = 12'b11110010_0_1;  // D18.7 (RD+)
      10'b1100101110: {data_o, k_char_o, valid_o} = 12'b11110011_0_1;  // D19.7 (RD-)
      10'b1100100001: {data_o, k_char_o, valid_o} = 12'b11110011_0_1;  // D19.7 (RD+)
      10'b0010110111: {data_o, k_char_o, valid_o} = 12'b11110100_0_1;  // D20.7 (RD-)
      10'b0010110001: {data_o, k_char_o, valid_o} = 12'b11110100_0_1;  // D20.7 (RD+)
      10'b1010101110: {data_o, k_char_o, valid_o} = 12'b11110101_0_1;  // D21.7 (RD-)
      10'b1010100001: {data_o, k_char_o, valid_o} = 12'b11110101_0_1;  // D21.7 (RD+)
      10'b0110101110: {data_o, k_char_o, valid_o} = 12'b11110110_0_1;  // D22.7 (RD-)
      10'b0110100001: {data_o, k_char_o, valid_o} = 12'b11110110_0_1;  // D22.7 (RD+)
      10'b1110100001: {data_o, k_char_o, valid_o} = 12'b11110111_0_1;  // D23.7 (RD+)
      10'b0001011110: {data_o, k_char_o, valid_o} = 12'b11110111_0_1;  // D23.7 (RD-)
      10'b1100110001: {data_o, k_char_o, valid_o} = 12'b11111000_0_1;  // D24.7 (RD+)
      10'b0011001110: {data_o, k_char_o, valid_o} = 12'b11111000_0_1;  // D24.7 (RD-)
      10'b1001101110: {data_o, k_char_o, valid_o} = 12'b11111001_0_1;  // D25.7 (RD-)
      10'b1001100001: {data_o, k_char_o, valid_o} = 12'b11111001_0_1;  // D25.7 (RD+)
      10'b0101101110: {data_o, k_char_o, valid_o} = 12'b11111010_0_1;  // D26.7 (RD-)
      10'b0101100001: {data_o, k_char_o, valid_o} = 12'b11111010_0_1;  // D26.7 (RD+)
      10'b1101100001: {data_o, k_char_o, valid_o} = 12'b11111011_0_1;  // D27.7 (RD+)
      10'b0010011110: {data_o, k_char_o, valid_o} = 12'b11111011_0_1;  // D27.7 (RD-)
      10'b0011101110: {data_o, k_char_o, valid_o} = 12'b11111100_0_1;  // D28.7 (RD-)
      10'b0011100001: {data_o, k_char_o, valid_o} = 12'b11111100_0_1;  // D28.7 (RD+)
      10'b1011100001: {data_o, k_char_o, valid_o} = 12'b11111101_0_1;  // D29.7 (RD+)
      10'b0100011110: {data_o, k_char_o, valid_o} = 12'b11111101_0_1;  // D29.7 (RD-)
      10'b0111100001: {data_o, k_char_o, valid_o} = 12'b11111110_0_1;  // D30.7 (RD+)
      10'b1000011110: {data_o, k_char_o, valid_o} = 12'b11111110_0_1;  // D30.7 (RD-)
      10'b1010110001: {data_o, k_char_o, valid_o} = 12'b11111111_0_1;  // D31.7 (RD+)
      10'b0101001110: {data_o, k_char_o, valid_o} = 12'b11111111_0_1;  // D31.7 (RD-)
      10'b0011110100: {data_o, k_char_o, valid_o} = 12'b00011100_1_1;  // K28.0 (RD+)
      10'b1100001011: {data_o, k_char_o, valid_o} = 12'b00011100_1_1;  // K28.0 (RD-)
      10'b0011111001: {data_o, k_char_o, valid_o} = 12'b00111100_1_1;  // K28.1 (RD+)
      10'b1100000110: {data_o, k_char_o, valid_o} = 12'b00111100_1_1;  // K28.1 (RD-)
      10'b0011110101: {data_o, k_char_o, valid_o} = 12'b01011100_1_1;  // K28.2 (RD+)
      10'b1100001010: {data_o, k_char_o, valid_o} = 12'b01011100_1_1;  // K28.2 (RD-)
      10'b0011110011: {data_o, k_char_o, valid_o} = 12'b01111100_1_1;  // K28.3 (RD+)
      10'b1100001100: {data_o, k_char_o, valid_o} = 12'b01111100_1_1;  // K28.3 (RD-)
      10'b0011110010: {data_o, k_char_o, valid_o} = 12'b10011100_1_1;  // K28.4 (RD+)
      10'b1100001101: {data_o, k_char_o, valid_o} = 12'b10011100_1_1;  // K28.4 (RD-)
      10'b0011111010: {data_o, k_char_o, valid_o} = 12'b10111100_1_1;  // K28.5 (RD+)
      10'b1100000101: {data_o, k_char_o, valid_o} = 12'b10111100_1_1;  // K28.5 (RD-)
      10'b0011110110: {data_o, k_char_o, valid_o} = 12'b11011100_1_1;  // K28.6 (RD+)
      10'b1100001001: {data_o, k_char_o, valid_o} = 12'b11011100_1_1;  // K28.6 (RD-)
      10'b0011111000: {data_o, k_char_o, valid_o} = 12'b11111100_1_1;  // K28.7 (RD+)
      10'b1100000111: {data_o, k_char_o, valid_o} = 12'b11111100_1_1;  // K28.7 (RD-)
      10'b1110101000: {data_o, k_char_o, valid_o} = 12'b11110111_1_1;  // K23.7 (RD+)
      10'b0001010111: {data_o, k_char_o, valid_o} = 12'b11110111_1_1;  // K23.7 (RD-)
      10'b1101101000: {data_o, k_char_o, valid_o} = 12'b11111011_1_1;  // K27.7 (RD+)
      10'b0010010111: {data_o, k_char_o, valid_o} = 12'b11111011_1_1;  // K27.7 (RD-)
      10'b1011101000: {data_o, k_char_o, valid_o} = 12'b11111101_1_1;  // K29.7 (RD+)
      10'b0100010111: {data_o, k_char_o, valid_o} = 12'b11111101_1_1;  // K29.7 (RD-)
      10'b0111101000: {data_o, k_char_o, valid_o} = 12'b11111110_1_1;  // K30.7 (RD+)
      10'b1000010111: {data_o, k_char_o, valid_o} = 12'b11111110_1_1;  // K30.7 (RD-)
      default:        {data_o, k_char_o, valid_o} = 12'b0000000000_0_0;  // ERROR
    endcase
  end

endmodule
